// Solutions for building from the waveforms
// circuit 1:
module top_module (
    input a,
    input b,
    output q );//

    assign q = a & b; // Fix me

endmodule

// circuit 2:

